** Profile: "Startup-trans"  [ c:\users\kesha\workspaces\odin\test\rotator\regulator\buck-boost\tps55165q1_12v_buck-boost_pspice_model\slvmca3a\tps55165-q1_pspice_trans\tps55165-q1_trans-pspicefiles\startup\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tps55165-q1_trans.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 14m 0 50n 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL2= 40
.OPTIONS ITL4= 60
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\Startup.net" 


.END
